library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity sign_ex is


    Port (	x  		: in std_logic_vector(15 downto 0);
				y			: out std_logic_vector(31 downto 0));
			  
		end sign_ex;
		
architecture Behavioral of sign_ex is
begin
	PROCESS(x)

		begin 
		if(x(15) = '1') then
			y(31) <= '1';
			y(30) <= '1';
			y(29) <= '1';
			y(28) <= '1';
			y(27) <= '1';
			y(26) <= '1';
			y(25) <= '1';
			y(24) <= '1';
			y(23) <= '1';
			y(22) <= '1';
			y(21) <= '1';
			y(20) <= '1';
			y(19) <= '1';
			y(18) <= '1';
			y(17) <= '1';
			y(16) <= '1';
			y(15) <= x(15);
			y(14) <= x(14);
			y(13) <= x(13);
			y(12) <= x(12);
			y(11) <= x(11);
			y(10) <= x(10);
			y(9) <= x(9);
			y(8) <= x(8);
			y(7) <= x(7);
			y(6) <= x(6);
			y(5) <= x(5);
			y(4) <= x(4);
			y(3) <= x(3);
			y(2) <= x(2);
			y(1) <= x(1);
			y(0) <= x(0);
		else
			y(31) <= '0';
			y(30) <= '0';
			y(29) <= '0';
			y(28) <= '0';
			y(27) <= '0';
			y(26) <= '0';
			y(25) <= '0';
			y(24) <= '0';
			y(23) <= '0';
			y(22) <= '0';
			y(21) <= '0';
			y(20) <= '0';
			y(19) <= '0';
			y(18) <= '0';
			y(17) <= '0';
			y(16) <= '0';
			y(15) <= x(15);
			y(14) <= x(14);
			y(13) <= x(13);
			y(12) <= x(12);
			y(11) <= x(11);
			y(10) <= x(10);
			y(9) <= x(9);
			y(8) <= x(8);
			y(7) <= x(7);
			y(6) <= x(6);
			y(5) <= x(5);
			y(4) <= x(4);
			y(3) <= x(3);
			y(2) <= x(2);
			y(1) <= x(1);
			y(0) <= x(0);
			
		end if;
	end process;

end Behavioral;